*******************************************************************************
*** CONTROL OPTIONS ***********************************************************
*******************************************************************************

*******************************************************************************
*** INCLUDES ******************************************************************
*******************************************************************************

*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.include 'deemb_kolding00_params.sp'

*******************************************************************************
*** SUBCIRCUITS ***************************************************************
*******************************************************************************

*******************************************************************************
*** CIRCUIT *******************************************************************
*******************************************************************************

P1 n1 GND port=1

RZcs1 n1 n1x 'Zc'
RZcg1 GND n1z 'Zc/2'
RZp1 n1x n1z 'Zp'
RZi1 n1x n1y 'Zi'
RZ11 n1z ncc 'Z1'
RZ31 n1y nc 'Z3'

RZf n1y n2y 'Zf'
RZ2 nc ncc 'Z2'

RZcs2 n2 n2x 'Zc'
RZcg2 GND2 n2z 'Zc/2'
RZp2 n2x n2z 'Zp'
RZi2 n2x n2y 'Zi'
RZ12 n2z ncc 'Z1'
RZ32 n2y nc 'Z3'

.model nmos S TSTONEFILE='deemb_dut.s2p'
Sdut n1y n2y nc mname=nmos

P2 n2 GND2 port=2

*******************************************************************************
*** ANALYSIS ******************************************************************
*******************************************************************************

.ac lin 100 1 300G
.lin sparcalc=1 format=touchstone filename=deemb_kolding00

*******************************************************************************
*** SAVED DATA ****************************************************************
*******************************************************************************

*******************************************************************************
*** HSPICE OPTIONS ************************************************************
*******************************************************************************

.option post nomod brief parhier=local

.end
