*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.param Zc=11
.param Zp=24e3
.param Z1=7
.param Z2=6
.param Z3=35e3
.param Zi=14
.param Zf=47e3
.param alpha=0.0

