*******************************************************************************
*** CONTROL OPTIONS ***********************************************************
*******************************************************************************

*******************************************************************************
*** INCLUDES ******************************************************************
*******************************************************************************

*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.include 'deemb_vandamme01_params.sp'

*******************************************************************************
*** SUBCIRCUITS ***************************************************************
*******************************************************************************

*******************************************************************************
*** CIRCUIT *******************************************************************
*******************************************************************************

P1 n1 GND port=1

RG1 n1 GND '1/G1'
RZ1 n1 n1x 'Z1'

RG3 n1x n2x '1/G3'
RZ3 nc GND 'Z3'

RG2 n2 GND '1/G2'
RZ2 n2 n2x 'Z2'

.model nmos S TSTONEFILE='deemb_dut.s2p'
Sdut n1x n2x nc mname=nmos

P2 n2 GND port=2

*******************************************************************************
*** ANALYSIS ******************************************************************
*******************************************************************************

.ac lin 100 1 300G
.lin sparcalc=1 format=touchstone filename=deemb_vandamme01

*******************************************************************************
*** SAVED DATA ****************************************************************
*******************************************************************************

*******************************************************************************
*** HSPICE OPTIONS ************************************************************
*******************************************************************************

.option post nomod brief parhier=local

.end
