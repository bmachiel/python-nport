*******************************************************************************
*** CONTROL OPTIONS ***********************************************************
*******************************************************************************

*******************************************************************************
*** INCLUDES ******************************************************************
*******************************************************************************

* from NCSU FreePDK45 [http://www.eda.ncsu.edu/wiki/FreePDK]
.include 'NMOS_VTG.inc'

*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.param W=4u
.param L=45n

.param Vg=0.7
.param Vd=0.7

*******************************************************************************
*** SUBCIRCUITS ***************************************************************
*******************************************************************************

*******************************************************************************
*** CIRCUIT *******************************************************************
*******************************************************************************

P1 n1x GND port=1 DC='Vg' RDC=0

M1 n2x n1x n3x n3x NMOS_VTG l='L' w='W' m=1

Rnul n3x GND 1e-5

P2 n2x GND port=2 DC='Vd' RDC=0

*******************************************************************************
*** ANALYSIS ******************************************************************
*******************************************************************************

.ac lin 100 1 300G
.lin sparcalc=1 format=touchstone filename=deemb_dut

*******************************************************************************
*** SAVED DATA ****************************************************************
*******************************************************************************

*******************************************************************************
*** HSPICE OPTIONS ************************************************************
*******************************************************************************

.option post nomod brief parhier=local

.end
