*******************************************************************************
*** CONTROL OPTIONS ***********************************************************
*******************************************************************************

*******************************************************************************
*** INCLUDES ******************************************************************
*******************************************************************************

*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.include 'deemb_twostep_params.sp'

*******************************************************************************
*** SUBCIRCUITS ***************************************************************
*******************************************************************************

*******************************************************************************
*** CIRCUIT *******************************************************************
*******************************************************************************

P1 n1 GND port=1

RY1 n1 GND '1/Y1'
RY2 n2 GND '1/Y2'
RY3 n1 n2 '1/Y3'

RZ1 n1 n1x 'Z1'
RZ2 n2 n2x 'Z2'
RZ3 nc GND 'Z3'

.model nmos S TSTONEFILE='deemb_dut.s2p'
Sdut n1x n2x nc mname=nmos

P2 n2 GND port=2

*******************************************************************************
*** ANALYSIS ******************************************************************
*******************************************************************************

.ac lin 100 1 300G
.lin sparcalc=1 format=touchstone filename=deemb_twostep

*******************************************************************************
*** SAVED DATA ****************************************************************
*******************************************************************************

*******************************************************************************
*** HSPICE OPTIONS ************************************************************
*******************************************************************************

.option post nomod brief parhier=local

.end
