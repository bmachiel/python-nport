* insert DUT into the S-parameters of the test fixture

*******************************************************************************
*** CONTROL OPTIONS ***********************************************************
*******************************************************************************

*******************************************************************************
*** INCLUDES ******************************************************************
*******************************************************************************

*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

*******************************************************************************
*** SUBCIRCUITS ***************************************************************
*******************************************************************************

*******************************************************************************
*** CIRCUIT *******************************************************************
*******************************************************************************

P1 n1 GND port=1

.model fixture S TSTONEFILE='deemb_mom_fixture.s4p'
Stestfixture n1 n2 n3 n4 GND mname=fixture

.model dut S TSTONEFILE='deemb_dut.s2p'
Sdut n3 n4 GND mname=dut

P2 n2 GND port=2

*******************************************************************************
*** ANALYSIS ******************************************************************
*******************************************************************************

.ac lin 100 1 110G
.lin sparcalc=1 format=touchstone filename=deemb_mom

*******************************************************************************
*** SAVED DATA ****************************************************************
*******************************************************************************

*******************************************************************************
*** HSPICE OPTIONS ************************************************************
*******************************************************************************

.option post nomod brief parhier=local

.end

