*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.param G1='1/24e3'
.param G2='1/35e3'
.param G3='1/47e3'
.param Z1=42
.param Z2=53
.param Z3=74

