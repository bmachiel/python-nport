*******************************************************************************
*** PARAMETERS ****************************************************************
*******************************************************************************

.param Y1='1/24e3'
.param Y2='1/35e3'
.param Y3='1/47e3'

.param Z1=42
.param Z2=53
.param Z3=74
